module csm #(
) (
    ports
);
    
endmodule